ENTITY nanoBlaze_tb IS
END nanoBlaze_tb;
